7 6 2 


