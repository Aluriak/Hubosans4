0 0 -1 -1 0 
0 1 -1 -1 0 
0 2 -1 -1 0 
0 3 -1 -1 0 
0 4 -1 -1 0 
0 5 -1 -1 0 
1 0 -1 -1 0 
1 1 -1 -1 0 
1 2 -1 -1 0 
1 3 -1 -1 0 
1 4 -1 -1 0 
1 5 -1 -1 0 
2 0 -1 -1 0 
2 1 -1 -1 0 
2 2 -1 -1 0 
2 3 -1 -1 0 
2 4 -1 -1 0 
2 5 -1 -1 0 
3 0 -1 -1 0 
3 1 -1 -1 0 
3 2 -1 -1 0 
3 3 -1 -1 0 
3 4 -1 -1 0 
3 5 -1 -1 0 
4 0 -1 -1 0 
4 1 -1 -1 0 
4 2 -1 -1 0 
4 3 -1 -1 0 
4 4 -1 -1 0 
4 5 -1 -1 0 
5 0 -1 -1 0 
5 1 -1 -1 0 
5 2 -1 -1 0 
5 3 -1 -1 0 
5 4 -1 -1 0 
5 5 -1 -1 0 
6 0 -1 -1 0 
6 1 -1 -1 0 
6 2 -1 -1 0 
6 3 -1 -1 0 
6 4 -1 -1 0 
6 5 -1 -1 0 
1 2 0 2 40 40 
0 0 33 0 1702195018 824210037 0 0 (null) 


